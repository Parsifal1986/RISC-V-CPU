module lsb (
  input wire clk,
  input wire rst,
  input wire rdy,
  input wire[7:0] mem_din,
  output wire[7:0] mem_dout,
  
)